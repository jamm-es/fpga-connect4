`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////
// generated with james's gen_sprite.py with arguments:
//     module_name: corner_border_check
//
//     image_file: sprites/corner_border_check.png
//     palette_file: palette.txt
//     canvas_width: 160
//     canvas_height: 120
//     x_offset: 0
//     y_offset: 0
//     x_tile: 1
//     y_tile: 1
//
//     inferred x bit length: 10
//     inferred y bit length: 10
//     inferred palette bit length: 4
//////////////////////////////////////////////////////////////////////////

module corner_border_check(clk, x, y, paletteIndex, valid);
    input wire clk;
    input wire[9:0] x;
    input wire[9:0] y;
    output reg[3:0] paletteIndex;
    output reg valid;

    reg [9:0] xOffset;
    reg [9:0] yOffset;
    reg [7:0] xSprite;
    reg [6:0] ySprite;
    reg inBounds;

    always @(posedge clk) begin
        xOffset = (x+0);
        yOffset = (y+0);
        xSprite = xOffset[7:0];
        ySprite = yOffset[6:0];
        inBounds = (xOffset >= 0 && xOffset < 160) && (yOffset >= 0 && yOffset < 120);

        case(ySprite)
            
            7'd0: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd1: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd2: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd3: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd4: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd5: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd6: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd7: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd8: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd9: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd10: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd11: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd12: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd13: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd14: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd15: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd16: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd17: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd18: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd19: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd20: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd21: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd22: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd23: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd24: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd25: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd26: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd27: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd28: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd29: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd30: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd31: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd32: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd33: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd34: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd35: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd36: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd37: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd38: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd39: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd40: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd41: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd42: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd43: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd44: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd45: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd46: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd47: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd48: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd49: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd50: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd51: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd52: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd53: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd54: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd55: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd56: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd57: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd58: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd59: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd60: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd61: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd62: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd63: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd64: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd65: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd66: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd67: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd68: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd69: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd70: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd71: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd72: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd73: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd74: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd75: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd76: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd77: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd78: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd79: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd80: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd81: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd82: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd83: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd84: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd85: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd86: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd87: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd88: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd89: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd90: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd91: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd92: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd93: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd94: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd95: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd96: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd97: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd98: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd99: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd100: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd101: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd102: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd103: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd104: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd105: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd106: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd107: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd108: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd109: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd110: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd111: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd112: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd113: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd114: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd115: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd2;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd116: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd117: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd118: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd15;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            
            7'd119: begin
               case(xSprite)
                    
                    8'd0: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd1: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd2: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd3: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd4: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd5: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd6: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd7: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd8: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd9: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd10: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd11: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd12: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd13: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd14: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd15: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd16: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd17: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd18: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd19: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd20: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd21: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd22: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd23: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd24: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd25: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd26: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd27: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd28: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd29: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd30: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd31: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd32: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd33: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd34: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd35: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd36: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd37: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd38: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd39: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd40: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd41: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd42: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd43: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd44: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd45: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd46: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd47: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd48: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd49: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd50: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd51: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd52: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd53: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd54: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd55: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd56: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd57: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd58: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd59: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd60: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd61: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd62: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd63: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd64: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd65: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd66: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd67: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd68: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd69: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd70: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd71: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd72: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd73: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd74: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd75: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd76: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd77: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd78: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd79: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd80: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd81: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd82: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd83: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd84: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd85: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd86: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd87: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd88: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd89: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd90: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd91: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd92: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd93: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd94: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd95: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd96: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd97: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd98: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd99: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd100: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd101: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd102: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd103: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd104: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd105: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd106: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd107: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd108: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd109: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd110: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd111: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd112: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd113: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd114: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd115: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd116: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd117: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd118: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd119: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd120: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd121: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd122: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd123: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd124: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd125: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd126: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd127: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd128: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd129: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd130: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd131: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd132: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd133: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd134: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd135: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd136: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd137: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd138: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd139: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd140: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd141: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd142: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd143: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd144: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd145: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd146: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd147: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd148: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd149: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd150: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd151: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd152: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd153: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd154: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd155: begin
                        paletteIndex = 4'd2;
                    end
                    
                    8'd156: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd157: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd158: begin
                        paletteIndex = 4'd12;
                    end
                    
                    8'd159: begin
                        paletteIndex = 4'd12;
                    end
                    

                    default: begin
                        paletteIndex = 4'bXXXX;
                    end
                endcase 
            end
            

            default: begin
                paletteIndex = 4'bXXXX;
            end
        endcase

        valid = inBounds && (paletteIndex != 4'd15);
    end


endmodule
